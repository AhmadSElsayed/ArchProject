LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


package Constants is
	constant OPCODE_NOP	: std_logic_vector(4 downto 0)	:= "00000";
	constant OPCODE_MOV	: std_logic_vector(4 downto 0)	:= "00001";
	constant OPCODE_ADD	: std_logic_vector(4 downto 0)	:= "00010";
	constant OPCODE_MUL	: std_logic_vector(4 downto 0)	:= "00011";
	constant OPCODE_SUB	: std_logic_vector(4 downto 0)	:= "00100";
	constant OPCODE_AND	: std_logic_vector(4 downto 0)	:= "00101";
	constant OPCODE_OR		: std_logic_vector(4 downto 0)	:= "00110";
	constant OPCODE_RLC	: std_logic_vector(4 downto 0)	:= "00111";
	constant OPCODE_RRC	: std_logic_vector(4 downto 0)	:= "01000";
	constant OPCODE_SHL	: std_logic_vector(4 downto 0)	:= "01001";
	constant OPCODE_SHR	: std_logic_vector(4 downto 0)	:= "01010";
	constant OPCODE_SETC	: std_logic_vector(4 downto 0)	:= "01011";
	constant OPCODE_CLRC	: std_logic_vector(4 downto 0)	:= "01100";
	constant OPCODE_PUSH	: std_logic_vector(4 downto 0)	:= "01101";
	constant OPCODE_POP	: std_logic_vector(4 downto 0)	:= "01110";
	constant OPCODE_OUT	: std_logic_vector(4 downto 0)	:= "01111";
	constant OPCODE_IN		: std_logic_vector(4 downto 0)	:= "10000";
	constant OPCODE_NOT	: std_logic_vector(4 downto 0)	:= "10001";
	constant OPCODE_NEG	: std_logic_vector(4 downto 0)	:= "10010";
	constant OPCODE_INC	: std_logic_vector(4 downto 0)	:= "10011";
	constant OPCODE_DEC	: std_logic_vector(4 downto 0)	:= "10100";
	constant OPCODE_JZ		: std_logic_vector(4 downto 0)	:= "10101";
	constant OPCODE_JN		: std_logic_vector(4 downto 0)	:= "10110";
	constant OPCODE_JC		: std_logic_vector(4 downto 0)	:= "10111";
	constant OPCODE_JMP	: std_logic_vector(4 downto 0)	:= "11000";
	constant OPCODE_CALL	: std_logic_vector(4 downto 0)	:= "11001";
	constant OPCODE_RET	: std_logic_vector(4 downto 0)	:= "11010";
	constant OPCODE_RTI	: std_logic_vector(4 downto 0)	:= "11011";
	constant OPCODE_LDM	: std_logic_vector(4 downto 0)	:= "11100";
	constant OPCODE_LDD	: std_logic_vector(4 downto 0)	:= "11101";
	constant OPCODE_STD	: std_logic_vector(4 downto 0)	:= "11110";
	constant OPCODE_ERROR	: std_logic_vector(4 downto 0)	:= "11111";
end package;